module io_interface(Address, IOR, IOW, Data);

/* Module Inputs */


endmodule
